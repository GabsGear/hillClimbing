* Circuit Name
M1 Vout VIN 0 0 N_1u l=1.5u w=3u
Rd VDD Vout 25000 
VDD VDD 0 5
vgss VIN N001 SINE(0 0.5 1) AC 1
VGS N001 0 1.5
.model NMOS NMOS
.model PMOS PMOS
.include cmosedu_models.txt
.meas gain FIND V(Vout)/V(Vin) AT 1
.tran 1s
.backanno
.end
