* Circuit Name
M1 Vout VIN 0 0 N_1u l=2.7935u w=21.8509u
Rd VDD Vout 45073.2
VDD VDD 0 5
vgss VIN N001 SINE(0 0.5 1) AC 1
VGS N001 0 1.11424
.model NMOS NMOS
.model PMOS PMOS
.include cmosedu_models.txt
.meas gain FIND V(Vout)/V(Vin) AT 1
.tran 1s
.backanno
.end
